interface intf(input clk,rst);
logic [3:0] in;
logic [1:0] s;
logic op;


endinterface