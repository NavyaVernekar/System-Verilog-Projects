`timescale 1ns / 1ps
interface intf(input sclk,rst);
logic cs;
logic mosi;
logic [15:0] data;

endinterface